	library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity T_FLIPFLOP_SOURCE is
   Port ( T,CLK,RES,TEMP : in  STD_LOGIC;
          Q,QB : out STD_LOGIC);
end T_FLIPFLOP_SOURCE;

architecture Behavioral of T_FLIPFLOP_SOURCE is

begin

PROCESS(T,CLK,RES)

VARIABLE TEMP:STD_LOGIC:='0';

BEGIN

IF(RES='1')THEN
TEMP:='0';
ELSIF(RISING_EDGE(CLK))THEN
IF(T='1')THEN
TEMP:= NOT TEMP;

END IF;
END IF;
Q<= NOT TEMP;
QB<= TEMP;

END PROCESS;
END BEHAVIORAL;